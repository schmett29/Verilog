// Verilog test fixture created from schematic C:\Users\luem\Desktop\lab03_dwe\lab03_dwe\PRELABTRIAL2.sch - Sun Sep 20 19:17:42 2015

`timescale 1ns / 1ps

module PRELABTRIAL2_PRELABTRIAL2_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   PRELABTRIAL2 UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
