// Verilog test fixture created from schematic C:\Users\bowditcw\lab06_dwe\nso_dwe.sch - Sun Oct 18 22:36:29 2015

`timescale 1ns / 1ps

module nso_dwe_nso_dwe_sch_tb();

// Inputs
   reg [6:0]S;
   reg L;
   reg R;
	reg Reset;

// Output
  wire [6:0]Sn;

// Bidirs

// Instantiate the UUT
   nso_dwe UUT (
		.S(S),
		.L(L), 
		.R(R), 
		.Reset(Reset),
		.Sn(Sn)
   );
// Initialize Inputs
   
       initial begin
		S = 7'b100000; #10;
		
		/*S0 = 1; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=0; Reset=0; #10;
		S0 = 1; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=1; Reset=0; #10;
		S0 = 1; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=0; Reset=0; #10;
		S0 = 1; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=1; Reset=0; #10;
		
		S0 = 0; S1 = 1; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=0; Reset=0; #10;
		S0 = 0; S1 = 1; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=1; Reset=0; #10;
		S0 = 0; S1 = 1; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=0; Reset=0; #10;
		S0 = 0; S1 = 1; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=1; Reset=0; #10;
		
		S0 = 0; S1 = 0; S2 = 1; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=0; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 1; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=0; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 1; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=1; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 1; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=1; Reset=0; #10;
		
		S0 = 0; S1 = 0; S2 = 0; S3 = 1; S4 = 0; S5 = 0; S6 = 0; L=0; R=0; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 1; S4 = 0; S5 = 0; S6 = 0; L=0; R=1; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 1; S4 = 0; S5 = 0; S6 = 0; L=1; R=0; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 1; S4 = 0; S5 = 0; S6 = 0; L=1; R=1; Reset=0; #10;
		
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 1; S5 = 0; S6 = 0; L=0; R=0; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 1; S5 = 0; S6 = 0; L=0; R=1; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 1; S5 = 0; S6 = 0; L=1; R=0; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 1; S5 = 0; S6 = 0; L=1; R=1; Reset=0; #10;
		
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 1; S6 = 0; L=0; R=0; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 1; S6 = 0; L=0; R=1; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 1; S6 = 0; L=1; R=0; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 1; S6 = 0; L=1; R=1; Reset=0; #10;
	
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 1; L=0; R=0; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 1; L=0; R=1; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 1; L=1; R=0; Reset=0; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 1; L=1; R=1; Reset=0; #10;
		
		
		S0 = 1; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=0; Reset=1; #10;
		S0 = 1; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=1; Reset=1; #10;
		S0 = 1; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=0; Reset=1; #10;
		S0 = 1; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=1; Reset=1; #10;
		
		S0 = 0; S1 = 1; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=0; Reset=1; #10;
		S0 = 0; S1 = 1; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=1; Reset=1; #10;
		S0 = 0; S1 = 1; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=0; Reset=1; #10;
		S0 = 0; S1 = 1; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=1; Reset=1; #10;
		
		S0 = 0; S1 = 0; S2 = 1; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=0; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 1; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=0; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 1; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=0; R=1; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 1; S3 = 0; S4 = 0; S5 = 0; S6 = 0; L=1; R=1; Reset=1; #10;
		
		S0 = 0; S1 = 0; S2 = 0; S3 = 1; S4 = 0; S5 = 0; S6 = 0; L=0; R=0; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 1; S4 = 0; S5 = 0; S6 = 0; L=0; R=1; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 1; S4 = 0; S5 = 0; S6 = 0; L=1; R=0; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 1; S4 = 0; S5 = 0; S6 = 0; L=1; R=1; Reset=1; #10;
		
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 1; S5 = 0; S6 = 0; L=0; R=0; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 1; S5 = 0; S6 = 0; L=0; R=1; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 1; S5 = 0; S6 = 0; L=1; R=0; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 1; S5 = 0; S6 = 0; L=1; R=1; Reset=1; #10;
		
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 1; S6 = 0; L=0; R=0; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 1; S6 = 0; L=0; R=1; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 1; S6 = 0; L=1; R=0; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 1; S6 = 0; L=1; R=1; Reset=1; #10;
	
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 1; L=0; R=0; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 1; L=0; R=1; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 1; L=1; R=0; Reset=1; #10;
		S0 = 0; S1 = 0; S2 = 0; S3 = 0; S4 = 0; S5 = 0; S6 = 1; L=1; R=1; Reset=1; #10;
		*/
		
   end
endmodule
